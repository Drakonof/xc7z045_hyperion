`define XILINX_PLATFORM