`timescale 1ns / 1ps

module sync_fifo_tb;






endmodule
